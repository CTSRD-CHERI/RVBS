// 2018, Alexandre Joannou, University of Cambridge

import DefaultValue :: *;
import RV_BasicTypes :: *;

import BID :: *;

///////////////////////////
// Interface to the CSRs //
////////////////////////////////////////////////////////////////////////////////

interface CSRs#(numeric type n);
  method ActionValue#(Bit#(n)) req (CSRReq#(n) r);
endinterface

typedef enum {RW, RS, RC} CSRReqType deriving (Eq, FShow);
typedef enum {ALL, NOREAD, NOWRITE} CSRReqEffects deriving (Eq, FShow);

typedef struct {
  Bit#(12) idx;
  Bit#(n) val;
  CSRReqType rType;
  CSRReqEffects rEffects;
} CSRReq#(numeric type n) deriving (FShow);

instance DefaultValue#(CSRReq#(n));
  function CSRReq#(n) defaultValue =
    CSRReq { idx: ?, val: ?, rType: RW, rEffects: ALL };
endinstance
function CSRReq#(n) rwCSRReq(Bit#(12) i, Bit#(n) v) =
  CSRReq { idx: i, val: v, rType: RW, rEffects: ALL };
function CSRReq#(n) rwCSRReqNoRead(Bit#(12) i, Bit#(n) v) =
  CSRReq { idx: i, val: v, rType: RW, rEffects: NOREAD };
function CSRReq#(n) rsCSRReq(Bit#(12) i, Bit#(n) v) =
  CSRReq { idx: i, val: v, rType: RS, rEffects: ALL };
function CSRReq#(n) rsCSRReqNoWrite(Bit#(12) i, Bit#(n) v) =
  CSRReq { idx: i, val: v, rType: RS, rEffects: NOWRITE };
function CSRReq#(n) rcCSRReq(Bit#(12) i, Bit#(n) v) =
  CSRReq { idx: i, val: v, rType: RC, rEffects: ALL };
function CSRReq#(n) rcCSRReqNoWrite(Bit#(12) i, Bit#(n) v) =
  CSRReq { idx: i, val: v, rType: RC, rEffects: NOWRITE };

//////////////////////////
// CSRs' implementation //
////////////////////////////////////////////////////////////////////////////////

function ActionValue#(Bit#(n)) readUpdateCSR(Reg#(csr_t) csr, CSRReq#(n) r)
provisos(Bits#(csr_t, n)) = actionvalue
  if (r.rEffects != NOWRITE) begin
    let newval = ?;
    case (r.rType)
      RW: newval = r.val;
      RS: newval = pack(csr) | r.val;
      RC: newval = pack(csr) & ~r.val;
    endcase
    csr <= unpack(newval);
    printTLogPlusArgs("CSRs", $format("overwriting 0x%0x with 0x%0x", pack(csr), newval));
  end
  return pack(csr);
endactionvalue;

function Bit#(2) xl_field(Integer xlen) = case (xlen)
  128: 2'b11; // 3
  64: 2'b10;  // 2
  32: 2'b01;  // 1
  default: 2'b00;
endcase;

////////////////////////
// machine level CSRs //
////////////////////////////////////////////////////////////////////////////////

typedef struct { Bit#(2) mxl; Bit#(TSub#(XLEN,28)) res; Bit#(26) extensions; }
  MISA deriving (Bits, FShow);
instance DefaultValue#(MISA);
  function MISA defaultValue() = MISA {
    `ifdef XLEN64
      mxl: 2'd2,
    `else
      mxl: 2'd1,
    `endif
    res: ?,
    extensions: 26'b00000000000000000100000000
  };
endinstance

typedef struct { Bit#(TSub#(XLEN,7)) bank; Bit#(7) offset; }
  MVENDORID deriving (Bits, FShow);
instance DefaultValue#(MVENDORID);
  function MVENDORID defaultValue() = MVENDORID {bank: 0, offset: 7'd0};
endinstance

typedef struct {
  Bool sd;
  `ifdef XLEN64 // MAX_XLEN > 32
  Bit#(TSub#(XLEN,37)) res4;
  Bit#(2) sxl;
  Bit#(2) uxl;
  Bit#(9) res3;
  `else // MAX_XLEN == 32
  Bit#(8) res3;
  `endif
  Bool tsr;
  Bool tw;
  Bool tvm;
  Bool mxr;
  Bool sum;
  Bool mprv;
  Bit#(2) xs;
  Bit#(2) fs;
  Bit#(2) mpp;
  Bit#(2) res2;
  Bool spp;
  Bool mpie;
  Bool res1;
  Bool spie;
  Bool upie;
  Bool mie;
  Bool res0;
  Bool sie;
  Bool uie;
} MSTATUS deriving (Bits, FShow);
instance DefaultValue#(MSTATUS);
  function MSTATUS defaultValue() = MSTATUS {
    sd: False,
    `ifdef XLEN64 // MAX_XLEN > 32
    res4: ?, sxl: xl_field(valueOf(XLEN)), uxl: xl_field(valueOf(XLEN)), res3: ?,
    `else // MAX_XLEN == 32
    res3: ?,
    `endif
    tsr: False, tw: False, tvm: False, mxr: False, sum: False, mprv: False,
    xs: 0, fs: 0, mpp: 0, res2: ?, spp: False,
    mpie: False, res1: ?, spie: False, upie: False,
    mie: False, res0: ?, sie: False, uie: False
  };
endinstance

//module [ArchStateDefModule#(n)] mkMCSRs(CSRs#(n))
module mkMCSRs(CSRs#(XLEN));

  // machine information registers
  //////////////////////////////////////////////////////////////////////////////
  Reg#(MVENDORID)  mvendorid <- mkReg(defaultValue); // mvendorid 12'hF11
  Reg#(Bit#(XLEN)) marchid   <- mkReg(0); // marchid 12'hF12
  Reg#(Bit#(XLEN)) mimpid    <- mkReg(0); // mimpid 12'hF13
  Reg#(Bit#(XLEN)) mhartid   <- mkReg(0); // mhartid 12'hF14

  // machine trap setup registers
  //////////////////////////////////////////////////////////////////////////////
  Reg#(MSTATUS)    mstatus <- mkReg(defaultValue); // mstatus 12'h300
  Reg#(MISA)       misa    <- mkReg(defaultValue); // misa 12'h301
  // medeleg 12'h302
  // mideleg 12'h303
  // mie 12'h304
  Reg#(Bit#(XLEN)) mtvec   <- mkReg(0); // mtvec 12'h305
  // mcounteren 12'h306

  // machine trap handling
  //////////////////////////////////////////////////////////////////////////////
  Reg#(Bit#(XLEN)) mscratch <- mkReg(0); // mscratch 12'h340
  // mepc 12'h341
  // mcause 12'h342
  // mtval 12'h343
  // mip 12'h344

  // machine protection and translation
  //////////////////////////////////////////////////////////////////////////////
  // pmpcfg0 12'h3A0
  // pmpcfg1 12'h3A1 (RV32 only)
  // pmpcfg2 12'h3A2
  // pmpcfg3 12'h3A3 (RV32 only)
  // pmpaddr0 12'h3B0
  // pmpaddr1 12'h3B1
  // ...
  // pmpaddr15 12'h3BF

  // machine CSR requests
  method ActionValue#(Bit#(XLEN)) req (CSRReq#(XLEN) r);
    Bit#(XLEN) ret = ?;
    case (r.idx) // TODO sort out individual behaviours for each CSR
      12'h300: ret <- readUpdateCSR(mstatus,r);
      12'h301: ret <- readUpdateCSR(misa,r);
      12'h305: ret <- readUpdateCSR(mtvec,r);
      12'h340: ret <- readUpdateCSR(mscratch,r);
      12'hF11: ret <- readUpdateCSR(mvendorid,r);
      12'hF12: ret <- readUpdateCSR(marchid,r);
      12'hF13: ret <- readUpdateCSR(mimpid,r);
      12'hF14: ret <- readUpdateCSR(mhartid,r);
      default: begin
        ret = ?;
        printLog($format("Machine CSR 0x%0x unimplemented - ", r.idx, fshow(r)));
      end
    endcase
    return ret;
  endmethod

endmodule

// user level CSRs
module [ArchStateDefModule#(XLEN)] mkUCSRs(CSRs#(XLEN));

  // user trap setup registers
  //////////////////////////////////////////////////////////////////////////////
  // ustatus 12'h000
  // uie 12'h004
  // utvec 12'h005

  // user trap handling
  //////////////////////////////////////////////////////////////////////////////
  // uscratch 12'h040
  // uepc 12'h041
  // ucause 12'h042
  // utval 12'h043
  // uip 12'h044

  // user counters/timers
  //////////////////////////////////////////////////////////////////////////////
  Reg#(Bit#(64)) cycle <- mkReg(0); // cycle 12'hC00 (and 12'hC80 in RV32)
  rule cycle_count;
    cycle <= cycle + 1;
  endrule
  // time 12'hC01 (and 12'hC81 in RV32)
  Reg#(Bit#(64)) instret <- mkCommittedInstCnt; // insret 12'hC02 (and 12'hC82 in RV32)
  // hpmcounter3 12'hC03 (and 12'hC83 in RV32)
  // hpmcounter4 12'hC04 (and 12'hC84 in RV32)
  // ...
  // hpmcounter31 12'hC1F (and 12'hC9F in RV32)

  method ActionValue#(Bit#(XLEN)) req (CSRReq#(XLEN) r);
    Bit#(XLEN) ret = ?;
    case (r.idx)
      12'hC00: ret = cycle[valueOf(XLEN)-1:0];
      12'hC02: ret = instret[valueOf(XLEN)-1:0];
      // RV32I only
      //'hC80: ret = cycle[63:32];
      //XXX hack for test suite
      12'hCC0: begin // test success
        $display("TEST SUCCESS");
        $finish(0);
      end
      12'hCC1: begin // test failure
        $display("TEST FAILURE");
        $finish(0);
      end
      default: begin
        ret = ?;
        printLog($format("User CSR 0x%0x unimplemented - ", r.idx, fshow(r)));
      end
    endcase
    return ret;
  endmethod

endmodule

module [ArchStateDefModule#(XLEN)] mkCSRs(CSRs#(XLEN));

  CSRs#(XLEN) uCSRs <- mkUCSRs;
  CSRs#(XLEN) mCSRs <- mkMCSRs;

  method ActionValue#(Bit#(XLEN)) req (CSRReq#(XLEN) r);
    printTLogPlusArgs("CSRs", $format("received ", fshow(r)));
    Bit#(XLEN) ret = ?;
    case (r.idx[9:8]) // lowest privilege level required for CSR access
      2'b00: ret <- uCSRs.req(r);
      2'b11: ret <- mCSRs.req(r);
      default: begin
        ret = ?;
        printLog($format("CSR 0x%0x unimplemented - ", r.idx, fshow(r)));
      end
    endcase
    return ret;
  endmethod

endmodule
