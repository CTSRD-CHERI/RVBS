// 2018, Alexandre Joannou, University of Cambridge

import RV_BasicTypes :: *;
export RV_BasicTypes :: *;

import RV_CSRs :: *;
export RV_CSRs :: *;

import RV_State :: *;
export RV_State :: *;

import RV_Mem :: *;
export RV_Mem :: *;

import RV_Trap :: *;
export RV_Trap :: *;
